// **************************************************
// ***************** Todo *************************** 
// **************************************************

// Delete parameters from read_data and write_data 

module Threshold
#(
    parameter 
        INPUT_FILE  = "input_picture.hex",  
        IMAGE_WIDTH = 768,                  
        IMAGE_HEIGHT = 512
    )
    (
        clk,                                                
        reset,                                  
                    
    );

    input clk;
    input reset;

endmodule 
